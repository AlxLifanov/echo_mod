/* Определение компонента Cping. На него ссылается класс echo.Server */

component echo.CPing // Название должно начинаться с большой буквы

endpoints {
    ping : echo.IPing  // Слева экземпляр интерфейса, справа его класс
}
