/* Определение компонента `ping`. На него ссылается класс echo.Server */

component echo.CPing

endpoints {
    ping : echo.IPing  // Название интерфейса, должно начинаться с большой буквы.
}
